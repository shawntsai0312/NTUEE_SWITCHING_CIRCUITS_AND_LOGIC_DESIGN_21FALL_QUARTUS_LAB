library verilog;
use verilog.vl_types.all;
entity AC4_vlg_vec_tst is
end AC4_vlg_vec_tst;
