library verilog;
use verilog.vl_types.all;
entity MU4_vlg_vec_tst is
end MU4_vlg_vec_tst;
