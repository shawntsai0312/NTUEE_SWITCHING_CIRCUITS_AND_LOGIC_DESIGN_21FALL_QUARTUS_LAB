library verilog;
use verilog.vl_types.all;
entity SD_vlg_vec_tst is
end SD_vlg_vec_tst;
