library verilog;
use verilog.vl_types.all;
entity FS4_vlg_vec_tst is
end FS4_vlg_vec_tst;
