library verilog;
use verilog.vl_types.all;
entity FA4_vlg_vec_tst is
end FA4_vlg_vec_tst;
