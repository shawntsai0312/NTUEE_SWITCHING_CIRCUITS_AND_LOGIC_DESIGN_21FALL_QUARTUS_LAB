library verilog;
use verilog.vl_types.all;
entity WSC_vlg_vec_tst is
end WSC_vlg_vec_tst;
